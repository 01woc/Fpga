module ecg_wave_gen (
    input clk,
    input reset,
    input [31:0] phase_acc,   // Đổi từ frequency thành phase_step
    output reg [23:0] ecg_wave // Sóng ECG đầu ra 24 bit
);

  
    reg [23:0] ecg_lut [0:1023]; // LUT chứa 1024 giá trị 24 bit

    // Khởi tạo LUT từ file
    initial begin
        $readmemh("D:/k242/Fgpa/fpga1.1/Fpga-main/Fpga-main/ecg_lut.dump", ecg_lut); // Nạp dữ liệu LUT từ file hex
    end

 

    // Tính địa chỉ LUT
    wire [9:0] lut_addr;
    assign lut_addr = phase_acc[31:22]; // Sử dụng 10 bit cao nhất của pha

    // Đọc giá trị sóng từ LUT
    always @(posedge clk) begin
        ecg_wave <= ecg_lut[lut_addr];
    end

endmodule
